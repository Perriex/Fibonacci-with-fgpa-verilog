module Controller();

endmodule