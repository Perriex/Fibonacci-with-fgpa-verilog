`timescale 1ns/1ns
module Datapath();

endmodule